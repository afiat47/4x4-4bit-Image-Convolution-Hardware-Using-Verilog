

`timescale 1ps / 1ps

module half_adder ( a ,b ,s ,c );

input a;
wire a;
input b;
wire b;
output s;
wire s;
output c;
wire c;			 


assign s = a ^ b;
assign c = a & b;



endmodule
